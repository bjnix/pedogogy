module part5(CLOCK_50,HEX7,HEX6,HEX5,HEX4,HEX3,HEX2,HEX1,HEX0);
	input CLOCK_50;
	output [6:0]HEX7,HEX6,HEX5,HEX4,HEX3,HEX2,HEX1,HEX0;
	
	reg [24:0] count;  //counter for clock
	
	//initial values for hex displays
	reg [2:0]d0= 3'b100; 
    reg [2:0]d1= 3'b011;
    reg [2:0]d2= 3'b010;
	reg	[2:0]d3= 3'b001;
	reg	[2:0]d4= 3'b000;
	reg	[2:0]d5= 3'b111;
	reg	[2:0]d6= 3'b110;
	reg	[2:0]d7= 3'b101;		
	
	always@ (posedge CLOCK_50)begin
			if (count == 0)begin
					d0=d0+1;
					d1=d1+1;
					d2=d2+1;
					d3=d3+1;
					d4=d4+1;
					d5=d5+1;
					d6=d6+1;
					d7=d7+1;
				end
				count=count+1; //counting action
			end
			
//outputs to displays
char_7seg s0(d0,HEX0);
char_7seg s1(d1,HEX1);
char_7seg s2(d2,HEX2);
char_7seg s3(d3,HEX3);
char_7seg s4(d4,HEX4);
char_7seg s5(d5,HEX5);
char_7seg s6(d6,HEX6);
char_7seg s7(d7,HEX7);


endmodule


//7-segment decoder
module char_7seg(C,Display);
	input[2:0]C;        
	output reg[6:0]Display; 
	
	
	always @(C)
		 case(C)
			3'b000 : Display =7'b1001000; //H
			3'b001 : Display =7'b0110000; //E
			3'b010 : Display =7'b1110001; //L
			3'b011 : Display =7'b1110001; //L
			3'b100 : Display =7'b0000001; //0
			default : Display =7'b1111111; //BLANK
		endcase	
endmodule
