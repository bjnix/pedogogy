module lab8(KEY,LEDR,LEDG,SW,HEX0,HEX1,HEX2,HEX3,HEX4,HEX5,HEX6,HEX7);
	input [17:0] SW;		//toggle switches
	input [1:0] KEY;
	output [6:0] HEX0;		//7-seg display 0 
	output [6:0] HEX1;		//"			  " 1
	output [6:0] HEX2; 		//"           " 2
	output [6:0] HEX3;		//"           " 3
	output [6:0] HEX4;		//"           " 4
	output [6:0] HEX5;		//"           " 5
	output [6:0] HEX6;		//"           " 6
	output [6:0] HEX7;		//"           " 7
	output [17:0] LEDR;		//red leds
	output [8:0]LEDG;

	
	wire [15:0] p0,p1,S;
	wire [7:0] A,B,C,D;
	reg [7:0] tmp0,tmp1;
	wire overflow;
	
	
	
	regi regiA (SW[15:8],KEY[1],KEY[0],(SW[17]&&SW[16]),A);
	regi regiB (SW[7:0],KEY[1],KEY[0],(SW[17]&&SW[16]),B);
	regi regiC (SW[15:8],KEY[1],KEY[0],(SW[17]&&(~SW[16])),C);
	regi regiD (SW[7:0],KEY[1],KEY[0],(SW[17]&&(~SW[16])),D);
	
	always@(SW[16],A,B,C,D) 
	begin
		if(SW[16])
			begin
				tmp0 = A;
				tmp1 = B;
			end
		else
			begin
				tmp0 = C;
				tmp1 = D;
			end
	end
	char_7seg h4(tmp1[3:0],HEX4);
	char_7seg h5(tmp1[7:4],HEX5);
	char_7seg h6(tmp0[3:0],HEX6);
	char_7seg h7(tmp0[7:4],HEX7);
	
	mult8 multab( A,B,p0 );
	mult8 multcd( C,D,p1 );
	addme addi( p0,p1,0,overflow,S );
	

	assign LEDG[8] = overflow; 
	// set output displays
	assign LEDR = {overflow,S};
	char_7seg h0(S[3:0],HEX0);
	char_7seg h1(S[7:4],HEX1);
	char_7seg h2(S[11:8],HEX2);
	char_7seg h3(S[15:12],HEX3);
	
endmodule 


module Oflow( D,Clk,Clr_n,Q );
	input Clk,Clr_n;
	input D;
	output reg Q;
	
	always@( negedge Clk, negedge Clr_n )
		begin
			if( !Clr_n )
				Q = 0;
			else
				Q = D;
		end
endmodule


module regi( D,Clk,Clr_n,enable,Q );
	input Clk,Clr_n,enable;
	input [7:0] D;
	output reg [7:0] Q;
	
	always@( negedge Clk, negedge Clr_n )
		begin
			if( !Clr_n )
				Q = 0;
			else if( Clr_n && enable )
				Q = D;
		end
endmodule


module full_adder ( A, B, C , M , Cout);
//A = input A
//B = input B
//C = input C
//M = result
//Cout = overflow bit 
	input A,B,C;
	output M,Cout;
	assign {Cout,M} = A + B + C;
		
endmodule
module char_7seg( C,Display );
	input[3:0]C;            //input code
	output reg[6:0]Display; //output 7-seg code
	
//assigns numbers to displays based on 4 bit input
	always@(C)
		case(C)
			4'b0000 : Display=7'b1000000; //0
			4'b0001 : Display=7'b1111001; //1
			4'b0010 : Display=7'b0100100; //2
			4'b0011 : Display=7'b0110000; //3
			4'b0100 : Display=7'b0011001; //4
			4'b0101 : Display=7'b0010010; //5
			4'b0110 : Display=7'b0000010; //6
			4'b0111 : Display=7'b1111000; //7
			4'b1000 : Display=7'b0000000; //8
			4'b1001 : Display=7'b0010000; //9
			4'b1010 : Display=7'b0001000; //A
			4'b1011 : Display=7'b0000011; //b
			4'b1100 : Display=7'b1000110; //c
			4'b1101 : Display=7'b0100001; //d
			4'b1110 : Display=7'b0000110; //E
			4'b1111 : Display=7'b0001110; //F
		endcase
	
endmodule

module addme(A,B,Cin,Cout,SUM);
	input [7:0] A,B;
	input Cin;
	output [7:0] SUM;
	output Cout;
	wire [7:0] M;
	wire [7:0] C;
	
	//------------------------- start add/subtract'n!
	//adder	
	full_adder fa0(A[0],B[0],   0,M[0],C[0]);
	full_adder fa1(A[1],B[1],C[0],M[1],C[1]);
	full_adder fa2(A[2],B[2],C[1],M[2],C[2]);
	full_adder fa3(A[3],B[3],C[2],M[3],C[3]);
	full_adder fa4(A[4],B[4],C[3],M[4],C[4]);
	full_adder fa5(A[5],B[5],C[4],M[5],C[5]);
	full_adder fa6(A[6],B[6],C[5],M[6],C[6]);
	full_adder fa7(A[7],B[7],C[6],M[7],C[7]);
	
	assign SUM = M;
	assign Cout = C[7];

endmodule
	
	
module mult8(A,B,P);
	input [7:0] A,B;
	output [15:0] P;
	wire [55:0] M,C;
//row0
	full_adder fa00(A[1]&B[0],A[0]&B[1],   0,M[0],C[0]);
	full_adder fa01(A[2]&B[0],A[1]&B[1],C[0],M[1],C[1]);
	full_adder fa02(A[3]&B[0],A[2]&B[1],C[1],M[2],C[2]);
	full_adder fa03(A[4]&B[0],A[3]&B[1],C[2],M[3],C[3]);
	full_adder fa04(A[5]&B[0],A[4]&B[1],C[3],M[4],C[4]);
	full_adder fa05(A[6]&B[0],A[5]&B[1],C[4],M[5],C[5]);
	full_adder fa06(A[7]&B[0],A[6]&B[1],C[5],M[6],C[6]);
	full_adder fa07(        0,A[7]&B[1],C[6],M[7],C[7]);
	//row1
	full_adder fa10(M[1],A[0]&B[2],0    ,M[ 8],C[ 8]);
	full_adder fa11(M[2],A[1]&B[2],C[ 8],M[ 9],C[ 9]);
	full_adder fa12(M[3],A[2]&B[2],C[ 9],M[10],C[10]);
	full_adder fa13(M[4],A[3]&B[2],C[10],M[11],C[11]);
	full_adder fa14(M[5],A[4]&B[2],C[11],M[12],C[12]);
	full_adder fa15(M[6],A[5]&B[2],C[12],M[13],C[13]);
	full_adder fa16(M[7],A[6]&B[2],C[13],M[14],C[14]);
	full_adder fa17(C[7],A[7]&B[2],C[14],M[15],C[15]);
	//row2
	full_adder fa20(M[ 9],A[0]&B[3],0    ,M[16],C[16]);
	full_adder fa21(M[10],A[1]&B[3],C[16],M[17],C[17]);
	full_adder fa22(M[11],A[2]&B[3],C[17],M[18],C[18]);
	full_adder fa23(M[12],A[3]&B[3],C[18],M[19],C[19]);
	full_adder fa24(M[13],A[4]&B[3],C[19],M[20],C[20]);
	full_adder fa25(M[14],A[5]&B[3],C[20],M[21],C[21]);
	full_adder fa26(M[15],A[6]&B[3],C[21],M[22],C[22]);
	full_adder fa27(C[15],A[7]&B[3],C[22],M[23],C[23]);
	//row3
	full_adder fa30(M[17],A[0]&B[4],0    ,M[24],C[24]);
	full_adder fa31(M[18],A[1]&B[4],C[24],M[25],C[25]);
	full_adder fa32(M[19],A[2]&B[4],C[25],M[26],C[26]);
	full_adder fa33(M[20],A[3]&B[4],C[26],M[27],C[27]);
	full_adder fa34(M[21],A[4]&B[4],C[27],M[28],C[28]);
	full_adder fa35(M[22],A[5]&B[4],C[28],M[29],C[29]);
	full_adder fa36(M[23],A[6]&B[4],C[29],M[30],C[30]);
	full_adder fa37(C[23],A[7]&B[4],C[30],M[31],C[31]);
	//row4
	full_adder fa40(M[25],A[0]&B[5],0    ,M[32],C[32]);
	full_adder fa41(M[26],A[1]&B[5],C[32],M[33],C[33]);
	full_adder fa42(M[27],A[2]&B[5],C[33],M[34],C[34]);
	full_adder fa43(M[28],A[3]&B[5],C[34],M[35],C[35]);
	full_adder fa44(M[29],A[4]&B[5],C[35],M[36],C[36]);
	full_adder fa45(M[30],A[5]&B[5],C[36],M[37],C[37]);
	full_adder fa46(M[31],A[6]&B[5],C[37],M[38],C[38]);
	full_adder fa47(C[31],A[7]&B[5],C[38],M[39],C[39]);
	//row5
	full_adder fa50(M[33],A[0]&B[6],0    ,M[40],C[40]);
	full_adder fa51(M[34],A[1]&B[6],C[40],M[41],C[41]);
	full_adder fa52(M[35],A[2]&B[6],C[41],M[42],C[42]);
	full_adder fa53(M[36],A[3]&B[6],C[42],M[43],C[43]);
	full_adder fa54(M[37],A[4]&B[6],C[43],M[44],C[44]);
	full_adder fa55(M[38],A[5]&B[6],C[44],M[45],C[45]);
	full_adder fa56(M[39],A[6]&B[6],C[45],M[46],C[46]);
	full_adder fa57(C[39],A[7]&B[6],C[46],M[47],C[47]);
	//row6
	full_adder fa60(M[41],A[0]&B[7],0    ,M[48],C[48]);
	full_adder fa61(M[42],A[1]&B[7],C[48],M[49],C[49]);
	full_adder fa62(M[43],A[2]&B[7],C[49],M[50],C[50]);
	full_adder fa63(M[44],A[3]&B[7],C[50],M[51],C[51]);
	full_adder fa64(M[45],A[4]&B[7],C[51],M[52],C[52]);
	full_adder fa65(M[46],A[5]&B[7],C[52],M[53],C[53]);
	full_adder fa66(M[47],A[6]&B[7],C[53],M[54],C[54]);
	full_adder fa67(C[47],A[7]&B[7],C[54],M[55],C[55]);
	
	assign P = {C[55],M[55],M[54],M[53],M[52],M[51],M[50],M[49],M[48],M[40],M[32],M[24],M[16],M[8],M[0],(A[0]&B[0])};
	
	
endmodule
	