//*/
module part2( Clk,D,Q );
	
	input Clk,D;
	output Q;
	
	wire R_g,S_g,Qa,Qb /*sythesis keep*/;
	
	assign R = ~D;
	assign S = D;
	
	nand( R_g,R,Clk );
	nand( S_g,S,Clk );
	nand( Qa,R_g,Qb );
	nand( Qb,S_g,Qa );

	assign Q = Qa;

endmodule